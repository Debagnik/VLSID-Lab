// Code your design here
module DFF(output Q,Qbar, input D,clk,rst);
  reg Q,Qbar;
  assign Qbar=!Q;
  always @(negedge clk) 
  begin
    if(rst==1)
      Q <= 0; 
    else 
      Q <= D; 
  end
endmodule 